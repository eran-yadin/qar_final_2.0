module label_generator (
    input sel,               // ����� �-SW[0] (���� ��� P1 �-P2)
    output [6:0] seg_P,      // ����� ��� �-Thousands (���� P)
    output reg [6:0] seg_num // ����� ��� �-Hundreds (1 �� 2)
);

    // ���� P �����
    assign seg_P = 7'b0001100; 

    always @(*) begin
        if (sel == 1'b0)
            seg_num = 7'b1111001; // ���� '1'
        else
            seg_num = 7'b0100100; // ���� '2'
    end

endmodule