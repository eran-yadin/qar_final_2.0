module pad_16_to_32_2 (
    input [15:0] data_in,   // ������ ������ (16 ���)
    output [31:0] data_out  // ������ �-BCD �� �-MUX (32 ���)
);

    // ����� ������� 16 ����� ��� ������ (����) �� �����
    assign data_out = {16'b0, data_in};

endmodule