module alu_32bit_2 (
    input [15:0] A,          // ���� ����� ����� 1
    input [15:0] B,          // ���� ��� ����� 2
    input [1:0]  op_select,  // ����� ����� (SW[9:8])
    output reg [31:0] result // ����� �-BCD
);

    // ����� ��� ������� ������ ����� �����
    reg [15:0] max_val;
    reg [15:0] min_val;

    always @(*) begin
        // ��� �������: ����� �� ����� ��� ����
        if (A >= B) begin
            max_val = A;
            min_val = B;
        end else begin
            max_val = B;
            min_val = A;
        end

        // ����� ������� ��� ������ ��������
        case (op_select)
            2'b00: result = {16'd0, (A + B)};          // ����� (���� ���)

            2'b01: result = {16'd0, (max_val - min_val)}; // �����: ���� ���� ���� ���

            2'b10: result = A*B;                     // ��� (���� ���)

            2'b11: begin                               // �����: ���� ���� ���� ���
                if (min_val != 0)
                    result = {16'd0, (max_val / min_val)};
                else
                    result = 32'hFFFFFFFF;            // ����� ����� ������ �-0
            end

            default: result = 32'd0;
        endcase
    end
endmodule