module demux_1to2_1bit (
    input data_in,   // ���� ����� (���� �-press �������)
    input sel,       // ��� ������ (���� SW0)
    output out0,     // ����� 0 (��� ����� A)
    output out1      // ����� 1 (��� ����� B)
);

    // ������ �����:
    // ������ ������� ����� �� �� sel ��� 0
    assign out0 = data_in & (~sel);
    
    // ������ ������ ����� �� �� sel ��� 1
    assign out1 = data_in & sel;

endmodule