module demux_1to2_16bit (
    input [15:0] data_in,    // ������ (16 ���)
    input sel,               // ��� ������ (0 �� 1)
    output reg [15:0] out0,  // ����� 0
    output reg [15:0] out1   // ����� 1
);

    always @(*) begin
        // ����� ����: ������� �������
        out0 = 16'd0;
        out1 = 16'd0;
        
        case (sel)
            1'b0: out0 = data_in; // ����� ����� ������ �������
            1'b1: out1 = data_in; // ����� ����� ������ ������
        endcase
    end
    
endmodule